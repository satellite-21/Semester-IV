`timescale 1ns / 1ps

module testCsa32Bit();
wire [31:0]sum;
wire cout;
reg [31:0]a;
reg [31:0]b;
carrySkip32 csa(a,b,sum,cout);
initial
    begin
    a=32'b00000000000000000000000000000000;b=32'b00000000000000000000000000000000;
    #100 a=32'b00000000000000000000000000000110;b=32'b00000000000000000000000000000100;
    #100 a=32'b00000000000000000000000000000010;b=32'b00000000000000000000000000000010;
    #100 a=32'b00000000000000000000000000000001;b=32'b00000000000000000000000000001000;
    end
initial #500 $finish;
endmodule